module auto_tune(CLOCK_50, left_audio_in,right_audio_in, left_audio_out, right_audio_out);


end module
